module calcdistance(in, out);
	input in;
	output out;
	wire [5:0] in;
	reg [11:0] out;
	
	always@(in)
	begin
		case (in)
			6'b000000:out <= 0;
			6'b000001:out <= 3300;
			6'b000010:out <= 1650;
			6'b000011:out <= 1100;
			6'b000100:out <= 825;
			6'b000101:out <= 660;
			6'b000110:out <= 550;
			6'b000111:out <= 471;
			6'b001000:out <= 412;
			6'b001001:out <= 366;
			6'b001010:out <= 330;
			6'b001011:out <= 300;
			6'b001100:out <= 275;
			6'b001101:out <= 253;
			6'b001110:out <= 235;
			6'b001111:out <= 220;
			6'b010000:out <= 206;
			6'b010001:out <= 194;
			6'b010010:out <= 183;
			6'b010011:out <= 173;
			6'b010100:out <= 165;
			6'b010101:out <= 157;
			6'b010110:out <= 150;
			6'b010111:out <= 143;
			6'b011000:out <= 137;
			6'b011001:out <= 132;
			6'b011010:out <= 126;
			6'b011011:out <= 122;
			6'b011100:out <= 117;
			6'b011101:out <= 113;
			6'b011110:out <= 110;
			6'b011111:out <= 106;
			6'b100000:out <= 103;
			6'b100001:out <= 100;
			6'b100010:out <= 97;
			6'b100011:out <= 94;
			6'b100100:out <= 91;
			6'b100101:out <= 89;
			6'b100110:out <= 86;
			6'b100111:out <= 84;
			6'b101000:out <= 82;
			6'b101001:out <= 80;
			6'b101010:out <= 78;
			6'b101011:out <= 76;
			6'b101100:out <= 75;
			6'b101101:out <= 73;
			6'b101110:out <= 71;
			6'b101111:out <= 70;
			6'b110000:out <= 68;
			6'b110001:out <= 67;
			6'b110010:out <= 66;
			6'b110011:out <= 64;
			6'b110100:out <= 63;
			6'b110101:out <= 62;
			6'b110110:out <= 61;
			6'b110111:out <= 60;
			6'b111000:out <= 58;
			6'b111001:out <= 57;
			6'b111010:out <= 56;
			6'b111011:out <= 55;
			6'b111100:out <= 55;
			6'b111101:out <= 54;
			6'b111110:out <= 53;
			6'b111111:out <= 52;
		endcase
	end
	
endmodule

