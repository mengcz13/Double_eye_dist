module formulacalc(sig, wf, f2sum, g2sum0, wg0, wfg0, fg0,
						g2sum1, wg1, wfg1, fg1,
						g2sum2, wg2, wfg2, fg2,
						g2sum3, wg3, wfg3, fg3,
						g2sum4, wg4, wfg4, fg4,
						g2sum5, wg5, wfg5, fg5,
						g2sum6, wg6, wfg6, fg6,
						g2sum7, wg7, wfg7, fg7,
						g2sum8, wg8, wfg8, fg8,
						g2sum9, wg9, wfg9, fg9,
						g2sum10, wg10, wfg10, fg10,
						g2sum11, wg11, wfg11, fg11,
						g2sum12, wg12, wfg12, fg12,
						g2sum13, wg13, wfg13, fg13,
						g2sum14, wg14, wfg14, fg14,
						g2sum15, wg15, wfg15, fg15,
						result);
	input sig;
	input wf, f2sum, g2sum0, wg0, wfg0, fg0;
	input g2sum1, wg1, wfg1, fg1;
	input g2sum2, wg2, wfg2, fg2;
	input g2sum3, wg3, wfg3, fg3; 
	input g2sum4, wg4, wfg4, fg4;
	input g2sum5, wg5, wfg5, fg5;
	input g2sum6, wg6, wfg6, fg6;
	input g2sum7, wg7, wfg7, fg7;
	input g2sum8, wg8, wfg8, fg8;
	input g2sum9, wg9, wfg9, fg9;
	input g2sum10, wg10, wfg10, fg10;
	input g2sum11, wg11, wfg11, fg11;
	input g2sum12, wg12, wfg12, fg12;
	input g2sum13, wg13, wfg13, fg13;
	input g2sum14, wg14, wfg14, fg14;
	input g2sum15, wg15, wfg15, fg15;
	
	wire sig;
	wire [13:0] wf;
	wire [13:0] f2sum;
	
	wire[55:0] g2sum0;
	wire[55:0] wg0;
	wire[55:0] wfg0;
	wire[55:0] fg0;
	wire[55:0] g2sum1;
	wire[55:0] wg1;
	wire[55:0] wfg1;
	wire[55:0] fg1;
	wire[55:0] g2sum2;
	wire[55:0] wg2;
	wire[55:0] wfg2;
	wire[55:0] fg2;
	wire[55:0] g2sum3;
	wire[55:0] wg3;
	wire[55:0] wfg3;
	wire[55:0] fg3;
	wire[55:0] g2sum4;
	wire[55:0] wg4;
	wire[55:0] wfg4;
	wire[55:0] fg4;
	wire[55:0] g2sum5;
	wire[55:0] wg5;
	wire[55:0] wfg5;
	wire[55:0] fg5;
	wire[55:0] g2sum6;
	wire[55:0] wg6;
	wire[55:0] wfg6;
	wire[55:0] fg6;
	wire[55:0] g2sum7;
	wire[55:0] wg7;
	wire[55:0] wfg7;
	wire[55:0] fg7;
	wire[55:0] g2sum8;
	wire[55:0] wg8;
	wire[55:0] wfg8;
	wire[55:0] fg8;
	wire[55:0] g2sum9;
	wire[55:0] wg9;
	wire[55:0] wfg9;
	wire[55:0] fg9;
	wire[55:0] g2sum10;
	wire[55:0] wg10;
	wire[55:0] wfg10;
	wire[55:0] fg10;
	wire[55:0] g2sum11;
	wire[55:0] wg11;
	wire[55:0] wfg11;
	wire[55:0] fg11;
	wire[55:0] g2sum12;
	wire[55:0] wg12;
	wire[55:0] wfg12;
	wire[55:0] fg12;
	wire[55:0] g2sum13;
	wire[55:0] wg13;
	wire[55:0] wfg13;
	wire[55:0] fg13;
	wire[55:0] g2sum14;
	wire[55:0] wg14;
	wire[55:0] wfg14;
	wire[55:0] fg14;
	wire[55:0] g2sum15;
	wire[55:0] wg15;
	wire[55:0] wfg15;
	wire[55:0] fg15;
	
	reg [1151:0] result; //18bit per block
	always@(posedge sig)
	begin;
		result[17:0] <= {0000, f2sum} + {0000, g2sum0[13:0]} + {000,wfg0[13:0], 0} - {0000, wf0[13:0]} - {0000, wg0[13:0]} - {000,fg0[13:0], 0};
		result[35:18] <= {0000, f2sum} + {0000, g2sum1[13:0]} + {000,wfg1[13:0], 0} - {0000, wf1[13:0]} - {0000, wg1[13:0]} - {000,fg1[13:0], 0};
		result[53:36] <= {0000, f2sum} + {0000, g2sum2[13:0]} + {000,wfg2[13:0], 0} - {0000, wf2[13:0]} - {0000, wg2[13:0]} - {000,fg2[13:0], 0};
		result[71:54] <= {0000, f2sum} + {0000, g2sum3[13:0]} + {000,wfg3[13:0], 0} - {0000, wf3[13:0]} - {0000, wg3[13:0]} - {000,fg3[13:0], 0};
		result[89:72] <= {0000, f2sum} + {0000, g2sum0[27:14]} + {000,wfg0[27:14], 0} - {0000, wf0[27:14]} - {0000, wg0[27:14]} - {000,fg0[27:14], 0};
		result[107:90] <= {0000, f2sum} + {0000, g2sum1[27:14]} + {000,wfg1[27:14], 0} - {0000, wf1[27:14]} - {0000, wg1[27:14]} - {000,fg1[27:14], 0};
		result[125:108] <= {0000, f2sum} + {0000, g2sum2[27:14]} + {000,wfg2[27:14], 0} - {0000, wf2[27:14]} - {0000, wg2[27:14]} - {000,fg2[27:14], 0};
		result[143:126] <= {0000, f2sum} + {0000, g2sum3[27:14]} + {000,wfg3[27:14], 0} - {0000, wf3[27:14]} - {0000, wg3[27:14]} - {000,fg3[27:14], 0};
		result[161:144] <= {0000, f2sum} + {0000, g2sum0[41:28]} + {000,wfg0[41:28], 0} - {0000, wf0[41:28]} - {0000, wg0[41:28]} - {000,fg0[41:28], 0};
		result[179:162] <= {0000, f2sum} + {0000, g2sum1[41:28]} + {000,wfg1[41:28], 0} - {0000, wf1[41:28]} - {0000, wg1[41:28]} - {000,fg1[41:28], 0};
		result[197:180] <= {0000, f2sum} + {0000, g2sum2[41:28]} + {000,wfg2[41:28], 0} - {0000, wf2[41:28]} - {0000, wg2[41:28]} - {000,fg2[41:28], 0};
		result[215:198] <= {0000, f2sum} + {0000, g2sum3[41:28]} + {000,wfg3[41:28], 0} - {0000, wf3[41:28]} - {0000, wg3[41:28]} - {000,fg3[41:28], 0};
		result[233:216] <= {0000, f2sum} + {0000, g2sum0[55:42]} + {000,wfg0[55:42], 0} - {0000, wf0[55:42]} - {0000, wg0[55:42]} - {000,fg0[55:42], 0};
		result[251:234] <= {0000, f2sum} + {0000, g2sum1[55:42]} + {000,wfg1[55:42], 0} - {0000, wf1[55:42]} - {0000, wg1[55:42]} - {000,fg1[55:42], 0};
		result[269:252] <= {0000, f2sum} + {0000, g2sum2[55:42]} + {000,wfg2[55:42], 0} - {0000, wf2[55:42]} - {0000, wg2[55:42]} - {000,fg2[55:42], 0};
		result[287:270] <= {0000, f2sum} + {0000, g2sum3[55:42]} + {000,wfg3[55:42], 0} - {0000, wf3[55:42]} - {0000, wg3[55:42]} - {000,fg3[55:42], 0};
		result[305:288] <= {0000, f2sum} + {0000, g2sum0[69:56]} + {000,wfg0[69:56], 0} - {0000, wf0[69:56]} - {0000, wg0[69:56]} - {000,fg0[69:56], 0};
		result[323:306] <= {0000, f2sum} + {0000, g2sum1[69:56]} + {000,wfg1[69:56], 0} - {0000, wf1[69:56]} - {0000, wg1[69:56]} - {000,fg1[69:56], 0};
		result[341:324] <= {0000, f2sum} + {0000, g2sum2[69:56]} + {000,wfg2[69:56], 0} - {0000, wf2[69:56]} - {0000, wg2[69:56]} - {000,fg2[69:56], 0};
		result[359:342] <= {0000, f2sum} + {0000, g2sum3[69:56]} + {000,wfg3[69:56], 0} - {0000, wf3[69:56]} - {0000, wg3[69:56]} - {000,fg3[69:56], 0};
		result[377:360] <= {0000, f2sum} + {0000, g2sum0[83:70]} + {000,wfg0[83:70], 0} - {0000, wf0[83:70]} - {0000, wg0[83:70]} - {000,fg0[83:70], 0};
		result[395:378] <= {0000, f2sum} + {0000, g2sum1[83:70]} + {000,wfg1[83:70], 0} - {0000, wf1[83:70]} - {0000, wg1[83:70]} - {000,fg1[83:70], 0};
		result[413:396] <= {0000, f2sum} + {0000, g2sum2[83:70]} + {000,wfg2[83:70], 0} - {0000, wf2[83:70]} - {0000, wg2[83:70]} - {000,fg2[83:70], 0};
		result[431:414] <= {0000, f2sum} + {0000, g2sum3[83:70]} + {000,wfg3[83:70], 0} - {0000, wf3[83:70]} - {0000, wg3[83:70]} - {000,fg3[83:70], 0};
		result[449:432] <= {0000, f2sum} + {0000, g2sum0[97:84]} + {000,wfg0[97:84], 0} - {0000, wf0[97:84]} - {0000, wg0[97:84]} - {000,fg0[97:84], 0};
		result[467:450] <= {0000, f2sum} + {0000, g2sum1[97:84]} + {000,wfg1[97:84], 0} - {0000, wf1[97:84]} - {0000, wg1[97:84]} - {000,fg1[97:84], 0};
		result[485:468] <= {0000, f2sum} + {0000, g2sum2[97:84]} + {000,wfg2[97:84], 0} - {0000, wf2[97:84]} - {0000, wg2[97:84]} - {000,fg2[97:84], 0};
		result[503:486] <= {0000, f2sum} + {0000, g2sum3[97:84]} + {000,wfg3[97:84], 0} - {0000, wf3[97:84]} - {0000, wg3[97:84]} - {000,fg3[97:84], 0};
		result[521:504] <= {0000, f2sum} + {0000, g2sum0[111:98]} + {000,wfg0[111:98], 0} - {0000, wf0[111:98]} - {0000, wg0[111:98]} - {000,fg0[111:98], 0};
		result[539:522] <= {0000, f2sum} + {0000, g2sum1[111:98]} + {000,wfg1[111:98], 0} - {0000, wf1[111:98]} - {0000, wg1[111:98]} - {000,fg1[111:98], 0};
		result[557:540] <= {0000, f2sum} + {0000, g2sum2[111:98]} + {000,wfg2[111:98], 0} - {0000, wf2[111:98]} - {0000, wg2[111:98]} - {000,fg2[111:98], 0};
		result[575:558] <= {0000, f2sum} + {0000, g2sum3[111:98]} + {000,wfg3[111:98], 0} - {0000, wf3[111:98]} - {0000, wg3[111:98]} - {000,fg3[111:98], 0};
		result[593:576] <= {0000, f2sum} + {0000, g2sum0[125:112]} + {000,wfg0[125:112], 0} - {0000, wf0[125:112]} - {0000, wg0[125:112]} - {000,fg0[125:112], 0};
		result[611:594] <= {0000, f2sum} + {0000, g2sum1[125:112]} + {000,wfg1[125:112], 0} - {0000, wf1[125:112]} - {0000, wg1[125:112]} - {000,fg1[125:112], 0};
		result[629:612] <= {0000, f2sum} + {0000, g2sum2[125:112]} + {000,wfg2[125:112], 0} - {0000, wf2[125:112]} - {0000, wg2[125:112]} - {000,fg2[125:112], 0};
		result[647:630] <= {0000, f2sum} + {0000, g2sum3[125:112]} + {000,wfg3[125:112], 0} - {0000, wf3[125:112]} - {0000, wg3[125:112]} - {000,fg3[125:112], 0};
		result[665:648] <= {0000, f2sum} + {0000, g2sum0[139:126]} + {000,wfg0[139:126], 0} - {0000, wf0[139:126]} - {0000, wg0[139:126]} - {000,fg0[139:126], 0};
		result[683:666] <= {0000, f2sum} + {0000, g2sum1[139:126]} + {000,wfg1[139:126], 0} - {0000, wf1[139:126]} - {0000, wg1[139:126]} - {000,fg1[139:126], 0};
		result[701:684] <= {0000, f2sum} + {0000, g2sum2[139:126]} + {000,wfg2[139:126], 0} - {0000, wf2[139:126]} - {0000, wg2[139:126]} - {000,fg2[139:126], 0};
		result[719:702] <= {0000, f2sum} + {0000, g2sum3[139:126]} + {000,wfg3[139:126], 0} - {0000, wf3[139:126]} - {0000, wg3[139:126]} - {000,fg3[139:126], 0};
		result[737:720] <= {0000, f2sum} + {0000, g2sum0[153:140]} + {000,wfg0[153:140], 0} - {0000, wf0[153:140]} - {0000, wg0[153:140]} - {000,fg0[153:140], 0};
		result[755:738] <= {0000, f2sum} + {0000, g2sum1[153:140]} + {000,wfg1[153:140], 0} - {0000, wf1[153:140]} - {0000, wg1[153:140]} - {000,fg1[153:140], 0};
		result[773:756] <= {0000, f2sum} + {0000, g2sum2[153:140]} + {000,wfg2[153:140], 0} - {0000, wf2[153:140]} - {0000, wg2[153:140]} - {000,fg2[153:140], 0};
		result[791:774] <= {0000, f2sum} + {0000, g2sum3[153:140]} + {000,wfg3[153:140], 0} - {0000, wf3[153:140]} - {0000, wg3[153:140]} - {000,fg3[153:140], 0};
		result[809:792] <= {0000, f2sum} + {0000, g2sum0[167:154]} + {000,wfg0[167:154], 0} - {0000, wf0[167:154]} - {0000, wg0[167:154]} - {000,fg0[167:154], 0};
		result[827:810] <= {0000, f2sum} + {0000, g2sum1[167:154]} + {000,wfg1[167:154], 0} - {0000, wf1[167:154]} - {0000, wg1[167:154]} - {000,fg1[167:154], 0};
		result[845:828] <= {0000, f2sum} + {0000, g2sum2[167:154]} + {000,wfg2[167:154], 0} - {0000, wf2[167:154]} - {0000, wg2[167:154]} - {000,fg2[167:154], 0};
		result[863:846] <= {0000, f2sum} + {0000, g2sum3[167:154]} + {000,wfg3[167:154], 0} - {0000, wf3[167:154]} - {0000, wg3[167:154]} - {000,fg3[167:154], 0};
		result[881:864] <= {0000, f2sum} + {0000, g2sum0[181:168]} + {000,wfg0[181:168], 0} - {0000, wf0[181:168]} - {0000, wg0[181:168]} - {000,fg0[181:168], 0};
		result[899:882] <= {0000, f2sum} + {0000, g2sum1[181:168]} + {000,wfg1[181:168], 0} - {0000, wf1[181:168]} - {0000, wg1[181:168]} - {000,fg1[181:168], 0};
		result[917:900] <= {0000, f2sum} + {0000, g2sum2[181:168]} + {000,wfg2[181:168], 0} - {0000, wf2[181:168]} - {0000, wg2[181:168]} - {000,fg2[181:168], 0};
		result[935:918] <= {0000, f2sum} + {0000, g2sum3[181:168]} + {000,wfg3[181:168], 0} - {0000, wf3[181:168]} - {0000, wg3[181:168]} - {000,fg3[181:168], 0};
		result[953:936] <= {0000, f2sum} + {0000, g2sum0[195:182]} + {000,wfg0[195:182], 0} - {0000, wf0[195:182]} - {0000, wg0[195:182]} - {000,fg0[195:182], 0};
		result[971:954] <= {0000, f2sum} + {0000, g2sum1[195:182]} + {000,wfg1[195:182], 0} - {0000, wf1[195:182]} - {0000, wg1[195:182]} - {000,fg1[195:182], 0};
		result[989:972] <= {0000, f2sum} + {0000, g2sum2[195:182]} + {000,wfg2[195:182], 0} - {0000, wf2[195:182]} - {0000, wg2[195:182]} - {000,fg2[195:182], 0};
		result[1007:990] <= {0000, f2sum} + {0000, g2sum3[195:182]} + {000,wfg3[195:182], 0} - {0000, wf3[195:182]} - {0000, wg3[195:182]} - {000,fg3[195:182], 0};
		result[1025:1008] <= {0000, f2sum} + {0000, g2sum0[209:196]} + {000,wfg0[209:196], 0} - {0000, wf0[209:196]} - {0000, wg0[209:196]} - {000,fg0[209:196], 0};
		result[1043:1026] <= {0000, f2sum} + {0000, g2sum1[209:196]} + {000,wfg1[209:196], 0} - {0000, wf1[209:196]} - {0000, wg1[209:196]} - {000,fg1[209:196], 0};
		result[1061:1044] <= {0000, f2sum} + {0000, g2sum2[209:196]} + {000,wfg2[209:196], 0} - {0000, wf2[209:196]} - {0000, wg2[209:196]} - {000,fg2[209:196], 0};
		result[1079:1062] <= {0000, f2sum} + {0000, g2sum3[209:196]} + {000,wfg3[209:196], 0} - {0000, wf3[209:196]} - {0000, wg3[209:196]} - {000,fg3[209:196], 0};
		result[1097:1080] <= {0000, f2sum} + {0000, g2sum0[223:210]} + {000,wfg0[223:210], 0} - {0000, wf0[223:210]} - {0000, wg0[223:210]} - {000,fg0[223:210], 0};
		result[1115:1098] <= {0000, f2sum} + {0000, g2sum1[223:210]} + {000,wfg1[223:210], 0} - {0000, wf1[223:210]} - {0000, wg1[223:210]} - {000,fg1[223:210], 0};
		result[1133:1116] <= {0000, f2sum} + {0000, g2sum2[223:210]} + {000,wfg2[223:210], 0} - {0000, wf2[223:210]} - {0000, wg2[223:210]} - {000,fg2[223:210], 0};
		result[1151:1134] <= {0000, f2sum} + {0000, g2sum3[223:210]} + {000,wfg3[223:210], 0} - {0000, wf3[223:210]} - {0000, wg3[223:210]} - {000,fg3[223:210], 0};
	end
endmodule