module calcdistance(in, out);
	input in;
	output out;
	wire [5:0] in;
	reg [11:0] out;
	
	always@(in)
	begin
		case (in)
			6'b000000:out <= 0;
			6'b000001:out <= 99;
			6'b000010:out <= 98;
			6'b000011:out <= 97;
			6'b000100:out <= 96;
			6'b000101:out <= 95;
			6'b000110:out <= 94;
			6'b000111:out <= 93;
			6'b001000:out <= 92;
			6'b001001:out <= 91;
			6'b001010:out <= 90;
			6'b001011:out <= 89;
			6'b001100:out <= 88;
			6'b001101:out <= 87;
			6'b001110:out <= 86;
			6'b001111:out <= 85;
			6'b010000:out <= 84;
			6'b010001:out <= 83;
			6'b010010:out <= 82;
			6'b010011:out <= 81;
			6'b010100:out <= 80;
			6'b010101:out <= 79;
			6'b010110:out <= 78;
			6'b010111:out <= 77;
			6'b011000:out <= 76;
			6'b011001:out <= 75;
			6'b011010:out <= 74;
			6'b011011:out <= 73;
			6'b011100:out <= 72;
			6'b011101:out <= 71;
			6'b011110:out <= 70;
			6'b011111:out <= 69;
			6'b100000:out <= 68;
			6'b100001:out <= 67;
			6'b100010:out <= 66;
			6'b100011:out <= 65;
			6'b100100:out <= 64;
			6'b100101:out <= 63;
			6'b100110:out <= 62;
			6'b100111:out <= 61;
			6'b101000:out <= 60;
			6'b101001:out <= 59;
			6'b101010:out <= 58;
			6'b101011:out <= 56;
			6'b101100:out <= 55;
			6'b101101:out <= 54;
			6'b101110:out <= 53;
			6'b101111:out <= 52;
			6'b110000:out <= 51;
			6'b110001:out <= 50;
			6'b110010:out <= 49;
			6'b110011:out <= 48;
			6'b110100:out <= 47;
			6'b110101:out <= 46;
			6'b110110:out <= 45;
			6'b110111:out <= 44;
			6'b111000:out <= 43;
			6'b111001:out <= 42;
			6'b111010:out <= 42;
			6'b111011:out <= 41;
			6'b111100:out <= 40;
			6'b111101:out <= 40;
			6'b111110:out <= 39;
			6'b111111:out <= 38;
		endcase
	end
	
endmodule

