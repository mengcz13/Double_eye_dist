module topcalc(data_in, clk, d);
	input clk;
	output d;
	
	calcfgs control {
		.clk(clk),
				
	};
	
	rightram right {
		.
	};
	
endmodule
