module binary2bcd(bn, Y_r);
input [3:0] bn;
output reg [6:0] Y_r;

always@(bn)
begin
case (bn)
4'b0000: Y_r = 7'b0111111; // 0
4'b0001: Y_r = 7'b0000110; // 1
4'b0010: Y_r = 7'b1011011; // 2
4'b0011: Y_r = 7'b1001111; // 3
4'b0100: Y_r = 7'b1100110; // 4
4'b0101: Y_r = 7'b1101101; // 5
4'b0110: Y_r = 7'b1111101; // 6
4'b0111: Y_r = 7'b0000111; // 7
4'b1000: Y_r = 7'b1111111; // 8
4'b1001: Y_r = 7'b1101111; // 9
4'b1010: Y_r = 7'b1110111; // A
4'b1011: Y_r = 7'b1111100; // b
4'b1100: Y_r = 7'b0111001; // c
4'b1101: Y_r = 7'b1011110; // d
4'b1110: Y_r = 7'b1111001; // E
4'b1111: Y_r = 7'b1110001; // F
default: Y_r = 7'b0000000;
endcase
end

endmodule