module coorcalc(x, y, z);
//坐标换算，输入图像的x与y坐标输出对应像素在RAM中对应的一维地址
//邹昊写
	input x, y;
	output z;
	wire [6:0] x;
	wire [3:0] y;
	reg [10:0] z;
	
	always@(x or y)
	begin
		case (y)
			4'b0000:z <= {4'b0000, x};
			4'b0001:z <= 11'b00001001111 + {4'b0000, x};
			4'b0010:z <= 11'b00010011110 + {4'b0000, x};
			4'b0011:z <= 11'b00011101101 + {4'b0000, x};
			4'b0100:z <= 11'b00100111100 + {4'b0000, x};
			4'b0101:z <= 11'b00110001011 + {4'b0000, x};
			4'b0110:z <= 11'b00111011010 + {4'b0000, x};
			4'b0111:z <= 11'b01000101001 + {4'b0000, x};
			4'b1000:z <= 11'b01001111000 + {4'b0000, x};
			4'b1001:z <= 11'b01011000111 + {4'b0000, x};
			4'b1010:z <= 11'b01100010110 + {4'b0000, x};
			4'b1011:z <= 11'b01101100101 + {4'b0000, x};
			4'b1100:z <= 11'b01110110100 + {4'b0000, x};
			4'b1101:z <= 11'b10000000011 + {4'b0000, x};
			4'b1110:z <= 11'b10001010010 + {4'b0000, x};
			4'b1111:z <= 11'b10010100001 + {4'b0000, x};
		endcase
	end
endmodule
